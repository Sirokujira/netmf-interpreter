/*
 * $Id: SimpleSample.cdl 1887 2012-09-14 07:26:36Z okuma-top $
 *
 * Simple �� Sample
 *
 *  +------------------------------------+           +----------------------+          +-------------+
 *  | mruby object                       |           |                      |          |             |
 *  |bridge=                             | sSample   |  tMrubyBridgesSample |  sSample |   tSample   |
 *  | TMrubyBridgesSampe("SimpleBridge") |==========>|     SimpleBridge     |----------|>  Sample    |
 *  |                                    |  �δؿ��� |                      |cCall eEnt|             |
 *  |                                    |           |                      |          |             |
 *  +------------------------------------+           +----------------------+          +-------------+
 *
 *�������˥��㵭��
 *
 *   sSample �� �ؿ����󥿥ե����������
 *              �����Ȥ�����Ƭʸ�� s ���ղä���
 * 
 *    �����˥��� sSample�ˤ� 2 �Ĥδؿ� sayHello �� howAreYou �����롣
 *    ���륿���� tSample ���󶡤��뵡ǽ�Ȥʤ�Τǡ�sSample �Ȥ���̾���ˤ�����
 *
 *�����륿���׵���
 *
 *   tMrubyBridgesSample �� �֥�å�����Υ��륿���� (MrubyBridgePlugin �ˤ������)
 *   tSample             �� �Ƥ���Υ��륿����
 *
 */

import( "cygwin_kernel.cdl" );

// �����˥��� sSample
signature sSample {
	ER  sayHello( [in]int32_t times );
	ER  howAreYou( [out,string(len)]char_t *buf, [in]int32_t len );
};

// ���륿���� tSample
celltype tSample {
	entry sSample eEnt;
};

// ���� Sample
cell tSample Sample
{
};

/*
 * �����˥���ץ饰���� MrubyBridgePlugin �θƤӽФ���
 *
 * MrubyBridgePlugin �ˤ��
 * ���֥�å��Υ��륿���� tMrubyBridgesSample ������� 
 *   gen/tmp_MrubyBridgePlugin_0.cdl ����������롣
 *   sSample ����ʬ�ϡ������˥���̾��
 * �����륿���ץ����� gen/tMrubyBridgesSample.c �ˡ�mruby �� 
 *   TMrubyBridgesSample ���饹��������ɤ���������롣
 */
generate( MrubyBridgePlugin, sSample, "" );

/*
 * �֥�å����������
 *
 * mruby ���顢TECS::tsSample ���饹�� Bridge �Ȥ��ƻ��Ȥ���롣
 *   ex) bridge = TECS::TsSample.new( "SimpleBridge" )
 *
 * cTECS �� signature�����ʤ�� sSample �δؿ�����TMrubyBridgesSample 
 * �Υ��󥹥��󥹥᥽�åɤȤ���������졢�ƤӽФ����Ȥ��Ǥ��롣
 *   ex) bridge.sayHello( 3 )
 */
cell nMruby::tsSample SimpleBridge {
  cTECS = Sample.eEnt;
};

// cell nMruby::tTECSInitializer VM_TECSInitializer;
cell nMruby::tMrubyProc VM {
  cInit = VM_TECSInitializer.eInitialize;
};

generate( C2TECSBridgePlugin, nPosix::sMain, "" );

cell nC2TECS::tnPosix_sMain Main {
	cCall = VM.eMain;
};
